`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// ECE369A - Computer Architecture
// Laboratory 1
// Module - ProgramCounter_tb.v
// Description - Test the 'ProgramCounter.v' module.
////////////////////////////////////////////////////////////////////////////////

module ProgramCounter_tb(); 

	reg [31:0] Address;
	reg Reset, Clk;

	wire [31:0] PCResult;

    ProgramCounter u0(
        .Address(Address), 
        .PCResult(PCResult), 
        .Reset(Reset), 
        .Clk(Clk)
    );

	initial begin
		Clk <= 1'b0;
		forever #10 Clk <= ~Clk;
	end

	initial begin
	
    /* Please fill in the implementation here... */
    
    /*Our testbench tests that when address is assigned some number, the Instruction
      (output) is the same. We also test that when rest is pressed, Instruction is
      set to 0*/
        @(posedge Clk);
        Reset <= 1'b1;
        @(posedge Clk);
        Reset <= 1'b0;
        @(posedge Clk);
        Address <= 1;
        @(posedge Clk);
        Address <= 10;
        @(posedge Clk);
        Reset <= 1;
	
	end

endmodule

